
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.subckt 1T1R_larger BL0 BL1 BE TE WL0 WL1 vddw gndw
N1 BE WL1 gndw gndw nhv
N0 TE WL0 gndw gndw nhv
X0 TE BE rram2 area_ox=0.1024 Tfilament_0=3.3e-9
P0 TE BL0 vddw vddw phv
P1 BE BL1 vddw vddw phv
.ends
